* CMOS Inverter – 0.5um – minArea Design
.include MOSFET_models_0p5_0p18-3.inc

* Power Supply
VDD  vdd  0  3.3

* Input source for DC sweep (will be overridden in .dc)
*Vin  in   0  3.3

* Load: RL + CL in series
Rload out n1 1k
Cload n1 0 0.5p
* MOSFETs
MNMOS out in 0 0 NMOS0P5 w=1.25u l=0.5u As=1.875p Ad=1.875p ps=5.5u pd=5.5u
MPMOS out in vdd vdd PMOS0P5 w=1.25u l=0.5u As=1.875p Ad=1.875p ps=5.5u pd=5.5u

* DC Sweep
*.dc Vin 0 3.3 0.005

* Operating point (optional)
*.op

* Transient input (enable during transient test)
Vin in 0 pulse(0 3.3 0 1p 1p 5n)

.tran 0.2n 10n
* Delay measurements (use only for transient)
.measure tpHL TRIG V(in) VAL=1.65 RISE=1  TARG V(out) VAL=1.65 FALL=1
.measure tpLH TRIG V(in) VAL=1.65 FALL=1  TARG V(out) VAL=1.65 RISE=1

.end
