* CMOS Inverter – 0.18um – Matched Design
.include MOSFET_models_0p5_0p18-3.inc

* Power Supply
VDD  vdd  0  1.8

* Input source for DC sweep (will be overridden in .dc)
*Vin  in   0  1.8

* Load: RL + CL in series
Rload out n1 1k
Cload n1 0 0.2p

* MOSFETs
MNMOS out in 0 0 NMOS0P18 w=0.9u l=0.18u As=0.486p Ad=0.486p ps=2.88u pd=2.88u
MPMOS out in vdd vdd PMOS0P18 w=4.05u l=0.18u As=2.187p Ad=2.187p ps=9.18u pd=9.18u

* DC Sweep
*.dc Vin 0 1.8 0.005

* Operating point (optional)
*.op

* Transient input (enable during transient test)
Vin in 0 pulse(0 1.8 0.2n 0.2n 0.2n 5n)

.tran 0.2n 10n
* Delay measurements (use only for transient)
*.measure tpHL TRIG V(in) VAL=0.9 RISE=1  TARG V(out) VAL=0.9 FALL=1
*.measure tpLH TRIG V(in) VAL=0.9 FALL=1  TARG V(out) VAL=0.9 RISE=1
* -------- Average Power Measurement Using INTEG ---------

* instantaneous power = V(VDD) * I(Vdd)
.measure TRAN P_integral INTEG ( V(VDD)*I(Vdd) ) FROM=0 TO=10n

* average power = integral / time window
.measure TRAN P_avg PARAM='P_integral / (10n - 0)'

.end
